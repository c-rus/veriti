--------------------------------------------------------------------------------
--! Project: veriti
--! Author: Chase Ruskin
--! Created: 2021-10-17
--! Package: veriti
--! Details:
--!     Low-level functions interacting between raw data layer and hardware 
--!     description for testbenches.
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library std;
use std.textio.all;

library work;
use work.casting;

package veriti is

    -- PUBLIC API

    --! Outputs a 50% duty cycle clock 'clk' with a period of 'period' that
    --! is continuously driven until 'halt' is set to 'true'. 
    procedure spin_clock(signal clk: out std_logic; period: time; signal halt: boolean);

    --! Asynchronously applies the reset (active-high) and then synchronously
    --! de-asserts the reset after 'cycles' clock cycles generated by 'clk'.
    --!
    --! The reset will not be applied if 'cycles' is set to 0. The reset will
    --! de-assert on the falling edge of the 'cycles' count clock cycle.
    procedure reset_system(signal clk: std_logic; signal rst: out std_logic; cycles: natural);

    --! Drive a logic vector signal in the testbench with a value from the file's row.
    procedure drive(variable row: inout line; signal vec: out std_logic_vector);

    --! Drive a logic vector signal in the testbench with a value from the file's row.
    procedure drive(variable row: inout line; signal wire: out std_logic);

    --! Read a logic vector variable's value form the file's row.
    procedure load(variable row: inout line; variable ideal: out std_logic_vector);

    --! Read a logic variable's value form the file's row.
    procedure load(variable row: inout line; variable ideal: out std_logic);

    --! Awaits the flag to be asserted or until delay time is up. Returns
    --! 'true' when the flag was asserted before the timeout and 'false' if
    --! the timeout was reached before the flag was raised.
    --!
    --! Sets an infinite delay if 'cycles' is set to 0.
    procedure monitor(signal clk: std_logic; signal flag: std_logic; cycles: natural; variable timeout: out boolean);

    --! Write a vector signal's value to the file's row.
    procedure store(variable row: inout line; vec: in std_logic_vector);
    
    --! Sets halt to 'true', prints a message to the console, and enters an
    --! infinite wait statement to signal that the simulation is complete.
    procedure complete(signal halt: out boolean);

    --! Enters infinite wait if the 'halt' signal is enabled.
    procedure check(halt: in boolean);

    --- ASSERTION FUNCTIONS

    procedure assert_eq(received: std_logic_vector; expected: std_logic_vector; comment: string);
    procedure assert_eq(received: std_logic; expected: std_logic; comment: string);

    procedure assert_ne(received: std_logic_vector; expected: std_logic_vector; comment: string);
    procedure assert_ne(received: std_logic; expected: std_logic; comment: string);

    procedure assert_stability(signal clk: std_logic; signal cond: std_logic; signal vec: std_logic_vector; comment: string);

    -- LOGGING FUNCTIONS

    procedure log(level: severity_level; comment: string);

    procedure err(comment: string);

end package;


package body veriti is

    procedure complete(signal halt: out boolean) is
    begin
        report "Simulation complete";
        halt <= true;
        wait;
    end procedure;

    procedure check(halt: in boolean) is
    begin
        if halt = true then 
            wait;
        end if;
    end procedure;


    procedure spin_clock(signal clk: out std_logic; period: time; signal halt: boolean) is
        variable inner_clk : std_logic := '0';
    begin
        while halt = false loop
            clk <= inner_clk;
            wait for period/2;
            inner_clk := not inner_clk;
        end loop;
        wait;
    end procedure;


    procedure reset_system(signal clk: std_logic; signal rst: out std_logic; cycles: natural) is
    begin
        -- only apply the reset if the number of cycles to delay is greater than zero
        if cycles > 0 then
            rst <= '1';
            wait for 0 ns;
            for delay in 1 to cycles loop
                wait until rising_edge(clk);
            end loop;
            wait until falling_edge(clk);
        end if;
        rst <= '0';
        -- wait for 0 ns;
    end procedure;


    procedure monitor(signal clk: std_logic; signal flag: std_logic; cycles: natural; variable timeout: out boolean) is
        variable cycle_count : natural := 0;
    begin
        timeout := true;
        if cycles = 0 then
            wait until rising_edge(clk) and flag = '1';
            timeout := false;
        else
            while cycle_count < cycles loop
                if flag = '1' then
                    timeout := false;
                    exit;
                end if;
                wait until rising_edge(clk);
                cycle_count := cycle_count + 1;
            end loop;
        end if;
    end procedure;


    procedure drive(variable row: inout line; signal vec: out std_logic_vector) is
        variable word      : string(vec'range);
        variable temp      : std_logic_vector(vec'range);
        variable delimiter : character;
    begin
        if row'length > 0 then
            read(row, word);
            for ii in vec'range loop
                temp(ii) := casting.char_to_logic(word(ii));
            end loop;
            vec <= temp;
            -- ignore the delimiter
            read(row, delimiter);
            -- wait for 0 ns;
        end if;
    end procedure;


    procedure load(variable row: inout line; variable ideal: out std_logic_vector) is
        variable word      : string(ideal'range);
        variable delimiter : character;
    begin
        if row'length > 0 then
            read(row, word);
            for ii in ideal'range loop
                ideal(ii) := casting.char_to_logic(word(ii));
            end loop;
            -- ignore the delimiter
            read(row, delimiter);
        end if;
    end procedure;


    procedure drive(variable row: inout line; signal wire: out std_logic) is
        variable word      : character;
        variable delimiter : character;
    begin
        if row'length > 0 then
            read(row, word);
            wire <= casting.char_to_logic(word);
            -- ignore the delimiter
            read(row, delimiter);
            -- wait for 0 ns;
        end if;
    end procedure;

    --! Read a signle-bit variable's value form the file's row.
    procedure load(variable row: inout line; variable ideal: out std_logic) is
        variable word      : character;
        variable delimiter : character;
    begin
        if row'length > 0 then
            read(row, word);
            ideal := casting.char_to_logic(word);
            -- ignore the delimiter
            read(row, delimiter);
        end if;
    end procedure;


    procedure store(variable row: inout line; vec: in std_logic_vector) is
        variable str : string(vec'range);
        variable str_index : positive := 1;
        variable delimiter : character := ',';
    begin
        for ii in vec'range loop
            if vec(ii) = '1' then
                str(ii) := '1';
            elsif vec(ii) = '0' then
                str(ii) := '0';
            else
                str(ii) := '?';
            end if;
        end loop;
        write(row, str);
        write(row, delimiter);
    end procedure;

    
    procedure log(level: severity_level; comment: string) is 
    begin
        if level = note then
            report "[NOTE]: " & comment severity note;
        elsif level = warning then
            report "[WARNING]: " & comment severity warning;
        elsif level = error then
            report "[ERROR]: " & comment severity error;
        elsif level = failure then
            report "[FAILURE]: " & comment severity failure;
        else 
            report "[INFO]: " & comment;
        end if;
    end procedure;


    procedure err(comment: string) is
    begin
        assert false report "[ERROR]: " & comment severity error;
    end procedure;


    procedure info(comment: string) is
    begin
        report "[INFO]: " & comment;
    end procedure;


    procedure assert_eq(received: std_logic_vector; expected: std_logic_vector; comment: string) is
    begin
        assert received = expected report 
            "[ERROR]: " & comment & " - " &
            "received " & casting.logics_to_str(received) & " != " &
            "expected " & casting.logics_to_str(expected)
        severity error;
    end procedure;

    procedure assert_eq(received: std_logic; expected: std_logic; comment: string) is
    begin
        assert received = expected report 
            "[ERROR]: " & comment & " - " &
            "received " & casting.logic_to_str(received) & " != " &
            "expected " & casting.logic_to_str(expected)
        severity error;
    end procedure;


    procedure assert_ne(received: std_logic_vector; expected: std_logic_vector; comment: string) is
    begin
        assert received /= expected report 
            "[ERROR]: " & comment & " - " &
            "received " & casting.logics_to_str(received) & " == " &
            "expected " & casting.logics_to_str(expected)
        severity error;
    end procedure;

    procedure assert_ne(received: std_logic; expected: std_logic; comment: string) is
    begin
        assert received /= expected report 
            "[ERROR]: " & comment & " - " &
            "received " & casting.logic_to_str(received) & " == " &
            "expected " & casting.logic_to_str(expected)
        severity error;
    end procedure;


    procedure assert_stability(signal clk: std_logic; signal cond: std_logic; signal vec: std_logic_vector; comment: string) is
        variable vec_prev: std_logic_vector(vec'range);
    begin
        wait until rising_edge(cond);
        -- wait until rising_edge(cond);
        vec_prev := vec;
        while cond = '1' loop
            -- check if its been stable since the rising edge of done
            assert vec_prev = vec report 
                "[ERROR]: " & comment & " - " &
                "updated value " & casting.logics_to_str(vec) & " != " &
                "assumed stability " & casting.logics_to_str(vec_prev)
            severity error;

            wait until rising_edge(clk);
        end loop;
    end procedure;



end package body;